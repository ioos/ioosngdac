netcdf IOOS_Glider_NetCDF_v3.0-qartod {
dimensions:
	time = UNLIMITED ; // (0 currently)
	traj_strlen = 20 ;
variables:
	char trajectory(traj_strlen) ;
		trajectory:cf_role = "trajectory_id" ;
		trajectory:comment = "A trajectory is a single deployment of a glider and may span multiple data files." ;
		trajectory:long_name = "Trajectory/Deployment Name" ;
	double time(time) ;
		time:ancillary_variables = "time_qc" ;
		time:calendar = "gregorian" ;
		time:comment = "Measured or calculated time at each point in the time-series" ;
		time:long_name = "Time" ;
		time:observation_type = "measured" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01T00:00:00Z" ;
	double lat(time) ;
		lat:_FillValue = -999. ;
		lat:ancillary_variables = "qartod_location_flag lat_qc" ;
		lat:comment = "Interpolated latitude at each point in the time-series" ;
		lat:coordinate_reference_frame = "urn:ogc:crs:EPSG::4326" ;
		lat:long_name = "Latitude" ;
		lat:observation_type = "measured" ;
		lat:platform = "platform" ;
		lat:reference = "WGS84" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:valid_max = 90. ;
		lat:valid_min = -90. ;
	double lon(time) ;
		lon:_FillValue = -999. ;
		lon:ancillary_variables = "qartod_location_flag lon_qc" ;
		lon:comment = "Interpolated longitude at each point in the time-series." ;
		lon:coordinate_reference_frame = "urn:ogc:crs:EPSG::4326" ;
		lon:long_name = "Longitude" ;
		lon:observation_type = "measured" ;
		lon:platform = "platform" ;
		lon:reference = "WGS84" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:valid_max = 180. ;
		lon:valid_min = -180. ;
	double pressure(time) ;
		pressure:_FillValue = -999. ;
		pressure:accuracy = " " ;
		pressure:ancillary_variables = "qartod_monotonic_pressure_flag qartod_pressure_flat_line_flag qartod_pressure_gross_range_flag qartod_pressure_rate_of_change_flag qartod_pressure_spike_flag pressure_qc" ;
		pressure:comment = " " ;
		pressure:instrument = "instrument_ctd" ;
		pressure:long_name = "Pressure" ;
		pressure:observation_type = "measured" ;
		pressure:platform = "platform" ;
		pressure:positive = "down" ;
		pressure:precision = " " ;
		pressure:reference_datum = "sea-surface" ;
		pressure:resolution = " " ;
		pressure:standard_name = "sea_water_pressure" ;
		pressure:units = "dbar" ;
		pressure:valid_max = 2000 ;
		pressure:valid_min = 0 ;
	double depth(time) ;
		depth:_FillValue = -999. ;
		depth:accuracy = " " ;
		depth:ancillary_variables = "depth_qc" ;
		depth:comment = " " ;
		depth:instrument = "instrument_ctd" ;
		depth:long_name = "Depth" ;
		depth:observation_type = "calculated" ;
		depth:platform = "platform" ;
		depth:positive = "down" ;
		depth:precision = " " ;
		depth:reference_datum = "sea-surface" ;
		depth:resolution = " " ;
		depth:standard_name = "depth" ;
		depth:units = "m" ;
		depth:valid_max = 2000 ;
		depth:valid_min = 0 ;
	double temperature(time) ;
		temperature:_FillValue = -999. ;
		temperature:accuracy = " " ;
		temperature:ancillary_variables = "qartod_temperature_climatological_flag qartod_temperature_flat_line_flag qartod_temperature_gross_range_flag qartod_temperature_rate_of_change_flag qartod_temperature_spike_flag temperature_qc" ;
		temperature:instrument = "instrument_ctd" ;
		temperature:long_name = "Temperature" ;
		temperature:observation_type = "measured" ;
		temperature:platform = "platform" ;
		temperature:precision = " " ;
		temperature:resolution = " " ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:units = "Celsius" ;
		temperature:valid_max = 40. ;
		temperature:valid_min = -5. ;
	double conductivity(time) ;
		conductivity:_FillValue = -999. ;
		conductivity:accuracy = " " ;
		conductivity:ancillary_variables = "qartod_conductivity_climatological_flag qartod_conductivity_flat_line_flag qartod_conductivity_gross_range_flag qartod_conductivity_rate_of_change_flag qartod_conductivity_spike_flag conductivity_qc" ;
		conductivity:instrument = "instrument_ctd" ;
		conductivity:long_name = "Conductivity" ;
		conductivity:observation_type = "measured" ;
		conductivity:platform = "platform" ;
		conductivity:precision = " " ;
		conductivity:resolution = " " ;
		conductivity:standard_name = "sea_water_electrical_conductivity" ;
		conductivity:units = "S m-1" ;
		conductivity:valid_max = 10. ;
		conductivity:valid_min = 0. ;
	double salinity(time) ;
		salinity:_FillValue = -999. ;
		salinity:accuracy = " " ;
		salinity:ancillary_variables = "qartod_salinity_climatological_flag qartod_salinity_flat_line_flag qartod_salinity_rate_of_change_flag qartod_salinity_spike_flag salinity_qc" ;
		salinity:instrument = "instrument_ctd" ;
		salinity:long_name = "Salinity" ;
		salinity:observation_type = "calculated" ;
		salinity:platform = "platform" ;
		salinity:precision = " " ;
		salinity:resolution = " " ;
		salinity:standard_name = "sea_water_practical_salinity" ;
		salinity:units = 1 ;
		salinity:valid_max = 40. ;
		salinity:valid_min = 0. ;
	double density(time) ;
		density:_FillValue = -999. ;
		density:accuracy = " " ;
		density:ancillary_variables = "qartod_density_climatological_flag qartod_density_flat_line_flag qartod_density_rate_of_change_flag qartod_density_spike_flag density_qc" ;
		density:instrument = "instrument_ctd" ;
		density:long_name = "Density" ;
		density:observation_type = "calculated" ;
		density:platform = "platform" ;
		density:precision = " " ;
		density:resolution = " " ;
		density:standard_name = "sea_water_density" ;
		density:units = "kg m-3" ;
		density:valid_max = 1040. ;
		density:valid_min = 1015. ;
	int profile_id ;
		profile_id:_FillValue = -999 ;
		profile_id:comment = "Sequential profile number within the trajectory.  This value is unique in each file that is part of a single trajectory/deployment." ;
		profile_id:long_name = "Profile ID" ;
		profile_id:valid_max = 2147483647 ;
		profile_id:valid_min = 1 ;
	double profile_time ;
		profile_time:_FillValue = -999. ;
		profile_time:calendar = "gregorian" ;
		profile_time:comment = "Timestamp corresponding to the mid-point of the profile" ;
		profile_time:long_name = "Profile Center Time" ;
		profile_time:observation_type = "calculated" ;
		profile_time:platform = "platform" ;
		profile_time:standard_name = "time" ;
		profile_time:units = "seconds since 1970-01-01T00:00:00Z" ;
	double profile_lat ;
		profile_lat:_FillValue = -999. ;
		profile_lat:comment = "Value is interpolated to provide an estimate of the latitude at the mid-point of the profile" ;
		profile_lat:long_name = "Profile Center Latitude" ;
		profile_lat:observation_type = "calculated" ;
		profile_lat:platform = "platform" ;
		profile_lat:standard_name = "latitude" ;
		profile_lat:units = "degrees_north" ;
		profile_lat:valid_max = 90. ;
		profile_lat:valid_min = -90. ;
	double profile_lon ;
		profile_lon:_FillValue = -999. ;
		profile_lon:comment = "Value is interpolated to provide an estimate of the longitude at the mid-point of the profile" ;
		profile_lon:long_name = "Profile Center Longitude" ;
		profile_lon:observation_type = "calculated" ;
		profile_lon:platform = "platform" ;
		profile_lon:standard_name = "longitude" ;
		profile_lon:units = "degrees_east" ;
		profile_lon:valid_max = 180. ;
		profile_lon:valid_min = -180. ;
	double time_uv ;
		time_uv:_FillValue = -999. ;
		time_uv:calendar = "gregorian" ;
		time_uv:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		time_uv:long_name = "Depth-Averaged Time" ;
		time_uv:observation_type = "calculated" ;
		time_uv:standard_name = "time" ;
		time_uv:units = "seconds since 1970-01-01T00:00:00Z" ;
	double lat_uv ;
		lat_uv:_FillValue = -999. ;
		lat_uv:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		lat_uv:long_name = "Depth-Averaged Latitude" ;
		lat_uv:observation_type = "calculated" ;
		lat_uv:platform = "platform" ;
		lat_uv:standard_name = "latitude" ;
		lat_uv:units = "degrees_north" ;
		lat_uv:valid_max = 90. ;
		lat_uv:valid_min = -90. ;
	double lon_uv ;
		lon_uv:_FillValue = -999. ;
		lon_uv:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		lon_uv:long_name = "Depth-Averaged Longitude" ;
		lon_uv:observation_type = "calculated" ;
		lon_uv:platform = "platform" ;
		lon_uv:standard_name = "longitude" ;
		lon_uv:units = "degrees_east" ;
		lon_uv:valid_max = 180. ;
		lon_uv:valid_min = -180. ;
	double u ;
		u:_FillValue = -999. ;
		u:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		u:long_name = "Depth-Averaged Eastward Sea Water Velocity" ;
		u:observation_type = "calculated" ;
		u:platform = "platform" ;
		u:standard_name = "eastward_sea_water_velocity" ;
		u:units = "m s-1" ;
		u:valid_max = 10. ;
		u:valid_min = -10. ;
	double v ;
		v:_FillValue = -999. ;
		v:comment = "The depth-averaged current is an estimate of the net current measured while the glider is underwater.  The value is calculated over the entire underwater segment, which may consist of 1 or more dives." ;
		v:long_name = "Depth-Averaged Northward Sea Water Velocity" ;
		v:observation_type = "calculated" ;
		v:platform = "platform" ;
		v:standard_name = "northward_sea_water_velocity" ;
		v:units = "m s-1" ;
		v:valid_max = 10. ;
		v:valid_min = -10. ;
	int platform ;
		platform:_FillValue = -999 ;
		platform:comment = " " ;
		platform:id = " " ;
		platform:instrument = "instrument_ctd" ;
		platform:long_name = " " ;
		platform:type = "platform" ;
		platform:wmo_id = " " ;
	int instrument_ctd ;
		instrument_ctd:_FillValue = -999 ;
		instrument_ctd:calibration_date = " " ;
		instrument_ctd:calibration_report = " " ;
		instrument_ctd:comment = "pumped CTD" ;
		instrument_ctd:factory_calibrated = " " ;
		instrument_ctd:long_name = "Seabird Glider Payload CTD" ;
		instrument_ctd:make_model = "Seabird GPCTD" ;
		instrument_ctd:platform = "platform" ;
		instrument_ctd:serial_number = " " ;
		instrument_ctd:type = "platform" ;
	byte time_qc(time) ;
		time_qc:_FillValue = -127b ;
		time_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		time_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		time_qc:long_name = "time Quality Flag" ;
		time_qc:standard_name = "time status_flag" ;
		time_qc:valid_max = 9b ;
		time_qc:valid_min = 0b ;
	byte lat_qc(time) ;
		lat_qc:_FillValue = -127b ;
		lat_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		lat_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		lat_qc:long_name = "lat Quality Flag" ;
		lat_qc:standard_name = "latitude status_flag" ;
		lat_qc:valid_max = 9b ;
		lat_qc:valid_min = 0b ;
	byte lon_qc(time) ;
		lon_qc:_FillValue = -127b ;
		lon_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		lon_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		lon_qc:long_name = "lon Quality Flag" ;
		lon_qc:standard_name = "longitude status_flag" ;
		lon_qc:valid_max = 9b ;
		lon_qc:valid_min = 0b ;
	byte pressure_qc(time) ;
		pressure_qc:_FillValue = -127b ;
		pressure_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		pressure_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		pressure_qc:long_name = "pressure Quality Flag" ;
		pressure_qc:standard_name = "sea_water_pressure status_flag" ;
		pressure_qc:valid_max = 9b ;
		pressure_qc:valid_min = 0b ;
	byte depth_qc(time) ;
		depth_qc:_FillValue = -127b ;
		depth_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		depth_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		depth_qc:long_name = "depth Quality Flag" ;
		depth_qc:standard_name = "depth status_flag" ;
		depth_qc:valid_max = 9b ;
		depth_qc:valid_min = 0b ;
	byte temperature_qc(time) ;
		temperature_qc:_FillValue = -127b ;
		temperature_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		temperature_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		temperature_qc:long_name = "temperature Quality Flag" ;
		temperature_qc:standard_name = "sea_water_temperature status_flag" ;
		temperature_qc:valid_max = 9b ;
		temperature_qc:valid_min = 0b ;
	byte conductivity_qc(time) ;
		conductivity_qc:_FillValue = -127b ;
		conductivity_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		conductivity_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		conductivity_qc:long_name = "conductivity Quality Flag" ;
		conductivity_qc:standard_name = "sea_water_electrical_conductivity status_flag" ;
		conductivity_qc:valid_max = 9b ;
		conductivity_qc:valid_min = 0b ;
	byte salinity_qc(time) ;
		salinity_qc:_FillValue = -127b ;
		salinity_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		salinity_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		salinity_qc:long_name = "salinity Quality Flag" ;
		salinity_qc:standard_name = "sea_water_practical_salinity status_flag" ;
		salinity_qc:valid_max = 9b ;
		salinity_qc:valid_min = 0b ;
	byte density_qc(time) ;
		density_qc:_FillValue = -127b ;
		density_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		density_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		density_qc:long_name = "density Quality Flag" ;
		density_qc:standard_name = "sea_water_density status_flag" ;
		density_qc:valid_max = 9b ;
		density_qc:valid_min = 0b ;
	byte profile_time_qc ;
		profile_time_qc:_FillValue = -127b ;
		profile_time_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		profile_time_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		profile_time_qc:long_name = "profile_time Quality Flag" ;
		profile_time_qc:standard_name = "time status_flag" ;
		profile_time_qc:valid_max = 9b ;
		profile_time_qc:valid_min = 0b ;
	byte profile_lat_qc ;
		profile_lat_qc:_FillValue = -127b ;
		profile_lat_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		profile_lat_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		profile_lat_qc:long_name = "profile_lat Quality Flag" ;
		profile_lat_qc:standard_name = "latitude status_flag" ;
		profile_lat_qc:valid_max = 9b ;
		profile_lat_qc:valid_min = 0b ;
	byte profile_lon_qc ;
		profile_lon_qc:_FillValue = -127b ;
		profile_lon_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		profile_lon_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		profile_lon_qc:long_name = "profile_lon Quality Flag" ;
		profile_lon_qc:standard_name = "longitude status_flag" ;
		profile_lon_qc:valid_max = 9b ;
		profile_lon_qc:valid_min = 0b ;
	byte time_uv_qc ;
		time_uv_qc:_FillValue = -127b ;
		time_uv_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		time_uv_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		time_uv_qc:long_name = "time_uv Quality Flag" ;
		time_uv_qc:standard_name = "time status_flag" ;
		time_uv_qc:valid_max = 9b ;
		time_uv_qc:valid_min = 0b ;
	byte lat_uv_qc ;
		lat_uv_qc:_FillValue = -127b ;
		lat_uv_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		lat_uv_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		lat_uv_qc:long_name = "lat_uv Quality Flag" ;
		lat_uv_qc:standard_name = "latitude status_flag" ;
		lat_uv_qc:valid_max = 9b ;
		lat_uv_qc:valid_min = 0b ;
	byte lon_uv_qc ;
		lon_uv_qc:_FillValue = -127b ;
		lon_uv_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		lon_uv_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		lon_uv_qc:long_name = "lon_uv Quality Flag" ;
		lon_uv_qc:standard_name = "longitude status_flag" ;
		lon_uv_qc:valid_max = 9b ;
		lon_uv_qc:valid_min = 0b ;
	byte u_qc ;
		u_qc:_FillValue = -127b ;
		u_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		u_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		u_qc:long_name = "u Quality Flag" ;
		u_qc:standard_name = "eastward_sea_water_velocity status_flag" ;
		u_qc:valid_max = 9b ;
		u_qc:valid_min = 0b ;
	byte v_qc ;
		v_qc:_FillValue = -127b ;
		v_qc:flag_meanings = "no_qc_performed good_data probably_good_data bad_data_that_are_potentially_correctable bad_data value_changed not_used not_used interpolated_value missing_value" ;
		v_qc:flag_values = 0b, 1b, 2b, 3b, 4b, 5b, 6b, 7b, 8b, 9b ;
		v_qc:long_name = "v Quality Flag" ;
		v_qc:standard_name = "northward_sea_water_velocity status_flag" ;
		v_qc:valid_max = 9b ;
		v_qc:valid_min = 0b ;
    // QARTOD Variables
    // Note these are optional and can be provided by data providers if QARTOD is performed.
	byte qartod_conductivity_climatological_flag(time) ;
		qartod_conductivity_climatological_flag:_FillValue = 9b ;
		qartod_conductivity_climatological_flag:long_name = "QARTOD conductivity climatological test" ;
		qartod_conductivity_climatological_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_conductivity_climatological_flag:valid_min = 1b ;
		qartod_conductivity_climatological_flag:valid_max = 4b ;
		qartod_conductivity_climatological_flag:flag_values = 1b, 3b, 4b ;
		qartod_conductivity_climatological_flag:comment = "QARTOD conductivity climatological test" ;
		qartod_conductivity_climatological_flag:standard_name = "sea_water_electrical_conductivity status_flag" ;
	byte qartod_conductivity_flat_line_flag(time) ;
		qartod_conductivity_flat_line_flag:_FillValue = 9b ;
		qartod_conductivity_flat_line_flag:long_name = "QARTOD conductivity flat line test" ;
		qartod_conductivity_flat_line_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_conductivity_flat_line_flag:valid_min = 1b ;
		qartod_conductivity_flat_line_flag:valid_max = 4b ;
		qartod_conductivity_flat_line_flag:flag_values = 1b, 3b, 4b ;
		qartod_conductivity_flat_line_flag:comment = "QARTOD conductivity flat line test" ;
		qartod_conductivity_flat_line_flag:standard_name = "sea_water_electrical_conductivity status_flag" ;
	byte qartod_conductivity_gross_range_flag(time) ;
		qartod_conductivity_gross_range_flag:_FillValue = 9b ;
		qartod_conductivity_gross_range_flag:long_name = "QARTOD conductivity gross range test" ;
		qartod_conductivity_gross_range_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_conductivity_gross_range_flag:valid_min = 1b ;
		qartod_conductivity_gross_range_flag:valid_max = 4b ;
		qartod_conductivity_gross_range_flag:flag_values = 1b, 3b, 4b ;
		qartod_conductivity_gross_range_flag:comment = "QARTOD conductivity gross range test" ;
		qartod_conductivity_gross_range_flag:standard_name = "sea_water_electrical_conductivity status_flag" ;
	byte qartod_conductivity_rate_of_change_flag(time) ;
		qartod_conductivity_rate_of_change_flag:_FillValue = 9b ;
		qartod_conductivity_rate_of_change_flag:long_name = "QARTOD conductivity rate of change test" ;
		qartod_conductivity_rate_of_change_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_conductivity_rate_of_change_flag:valid_min = 1b ;
		qartod_conductivity_rate_of_change_flag:valid_max = 4b ;
		qartod_conductivity_rate_of_change_flag:flag_values = 1b, 3b, 4b ;
		qartod_conductivity_rate_of_change_flag:comment = "QARTOD conductivity rate of change test" ;
		qartod_conductivity_rate_of_change_flag:standard_name = "sea_water_electrical_conductivity status_flag" ;
	byte qartod_conductivity_spike_flag(time) ;
		qartod_conductivity_spike_flag:_FillValue = 9b ;
		qartod_conductivity_spike_flag:long_name = "QARTOD conductivity spike test" ;
		qartod_conductivity_spike_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_conductivity_spike_flag:valid_min = 1b ;
		qartod_conductivity_spike_flag:valid_max = 4b ;
		qartod_conductivity_spike_flag:flag_values = 1b, 3b, 4b ;
		qartod_conductivity_spike_flag:comment = "QARTOD conductivity spike test" ;
		qartod_conductivity_spike_flag:standard_name = "sea_water_electrical_conductivity status_flag" ;
	byte qartod_density_climatological_flag(time) ;
		qartod_density_climatological_flag:_FillValue = 9b ;
		qartod_density_climatological_flag:long_name = "QARTOD density climatology test" ;
		qartod_density_climatological_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_density_climatological_flag:valid_min = 1b ;
		qartod_density_climatological_flag:valid_max = 4b ;
		qartod_density_climatological_flag:flag_values = 1b, 3b, 4b ;
		qartod_density_climatological_flag:comment = "QARTOD density climatology test" ;
		qartod_density_climatological_flag:standard_name = "sea_water_density status_flag" ;
	byte qartod_density_flat_line_flag(time) ;
		qartod_density_flat_line_flag:_FillValue = 9b ;
		qartod_density_flat_line_flag:long_name = "QARTOD density flat line test" ;
		qartod_density_flat_line_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_density_flat_line_flag:valid_min = 1b ;
		qartod_density_flat_line_flag:valid_max = 4b ;
		qartod_density_flat_line_flag:flag_values = 1b, 3b, 4b ;
		qartod_density_flat_line_flag:comment = "QARTOD density flat line test" ;
		qartod_density_flat_line_flag:standard_name = "sea_water_density status_flag" ;
	byte qartod_density_rate_of_change_flag(time) ;
		qartod_density_rate_of_change_flag:_FillValue = 9b ;
		qartod_density_rate_of_change_flag:long_name = "QARTOD density rate of change test" ;
		qartod_density_rate_of_change_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_density_rate_of_change_flag:valid_min = 1b ;
		qartod_density_rate_of_change_flag:valid_max = 4b ;
		qartod_density_rate_of_change_flag:flag_values = 1b, 3b, 4b ;
		qartod_density_rate_of_change_flag:comment = "QARTOD density rate of change test" ;
		qartod_density_rate_of_change_flag:standard_name = "sea_water_density status_flag" ;
	byte qartod_density_spike_flag(time) ;
		qartod_density_spike_flag:_FillValue = 9b ;
		qartod_density_spike_flag:long_name = "QARTOD density spike test" ;
		qartod_density_spike_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_density_spike_flag:valid_min = 1b ;
		qartod_density_spike_flag:valid_max = 4b ;
		qartod_density_spike_flag:flag_values = 1b, 3b, 4b ;
		qartod_density_spike_flag:comment = "QARTOD density spike test" ;
		qartod_density_spike_flag:standard_name = "sea_water_density status_flag" ;
	byte qartod_location_flag ;
		qartod_location_flag:_FillValue = 9b ;
		qartod_location_flag:long_name = "QARTOD location test" ;
		qartod_location_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_location_flag:valid_min = 1b ;
		qartod_location_flag:valid_max = 4b ;
		qartod_location_flag:flag_values = 1b, 3b, 4b ;
		qartod_location_flag:comment = "QARTOD location test" ;
	byte qartod_monotonic_pressure_flag(time) ;
		qartod_monotonic_pressure_flag:_FillValue = 9b ;
		qartod_monotonic_pressure_flag:long_name = "QARTOD monotonic pressure test" ;
		qartod_monotonic_pressure_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_monotonic_pressure_flag:valid_min = 1b ;
		qartod_monotonic_pressure_flag:valid_max = 4b ;
		qartod_monotonic_pressure_flag:flag_values = 1b, 3b, 4b ;
		qartod_monotonic_pressure_flag:comment = "QARTOD monotonic pressure test" ;
		qartod_monotonic_pressure_flag:standard_name = "sea_water_pressure status_flag" ;
	byte qartod_pressure_flat_line_flag(time) ;
		qartod_pressure_flat_line_flag:_FillValue = 9b ;
		qartod_pressure_flat_line_flag:long_name = "QARTOD pressure flat line test" ;
		qartod_pressure_flat_line_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_pressure_flat_line_flag:valid_min = 1b ;
		qartod_pressure_flat_line_flag:valid_max = 4b ;
		qartod_pressure_flat_line_flag:flag_values = 1b, 3b, 4b ;
		qartod_pressure_flat_line_flag:comment = "QARTOD pressure flat line test" ;
		qartod_pressure_flat_line_flag:standard_name = "sea_water_pressure status_flag" ;
	byte qartod_pressure_gross_range_flag(time) ;
		qartod_pressure_gross_range_flag:_FillValue = 9b ;
		qartod_pressure_gross_range_flag:long_name = "QARTOD pressure gross range test" ;
		qartod_pressure_gross_range_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_pressure_gross_range_flag:valid_min = 1b ;
		qartod_pressure_gross_range_flag:valid_max = 4b ;
		qartod_pressure_gross_range_flag:flag_values = 1b, 3b, 4b ;
		qartod_pressure_gross_range_flag:comment = "QARTOD pressure gross range test" ;
		qartod_pressure_gross_range_flag:standard_name = "sea_water_pressure status_flag" ;
	byte qartod_pressure_rate_of_change_flag(time) ;
		qartod_pressure_rate_of_change_flag:_FillValue = 9b ;
		qartod_pressure_rate_of_change_flag:long_name = "QARTOD pressure rate of change" ;
		qartod_pressure_rate_of_change_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_pressure_rate_of_change_flag:valid_min = 1b ;
		qartod_pressure_rate_of_change_flag:valid_max = 4b ;
		qartod_pressure_rate_of_change_flag:flag_values = 1b, 3b, 4b ;
		qartod_pressure_rate_of_change_flag:comment = "QARTOD pressure rate of change test" ;
		qartod_pressure_rate_of_change_flag:standard_name = "sea_water_pressure status_flag" ;
	byte qartod_pressure_spike_flag(time) ;
		qartod_pressure_spike_flag:_FillValue = 9b ;
		qartod_pressure_spike_flag:long_name = "QARTOD pressure spike test" ;
		qartod_pressure_spike_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_pressure_spike_flag:valid_min = 1b ;
		qartod_pressure_spike_flag:valid_max = 4b ;
		qartod_pressure_spike_flag:flag_values = 1b, 3b, 4b ;
		qartod_pressure_spike_flag:comment = "QARTOD pressure spike test" ;
		qartod_pressure_spike_flag:standard_name = "sea_water_pressure status_flag" ;
	byte qartod_salinity_climatological_flag(time) ;
		qartod_salinity_climatological_flag:_FillValue = 9b ;
		qartod_salinity_climatological_flag:long_name = "QARTOD salinity climatological test" ;
		qartod_salinity_climatological_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_salinity_climatological_flag:valid_min = 1b ;
		qartod_salinity_climatological_flag:valid_max = 4b ;
		qartod_salinity_climatological_flag:flag_values = 1b, 3b, 4b ;
		qartod_salinity_climatological_flag:comment = "QARTOD salinity climatological test" ;
		qartod_salinity_climatological_flag:standard_name = "sea_water_salinity status_flag" ;
	byte qartod_salinity_flat_line_flag(time) ;
		qartod_salinity_flat_line_flag:_FillValue = 9b ;
		qartod_salinity_flat_line_flag:long_name = "QARTOD salinity flat line test" ;
		qartod_salinity_flat_line_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_salinity_flat_line_flag:valid_min = 1b ;
		qartod_salinity_flat_line_flag:valid_max = 4b ;
		qartod_salinity_flat_line_flag:flag_values = 1b, 3b, 4b ;
		qartod_salinity_flat_line_flag:comment = "QARTOD salinity flat line test" ;
		qartod_salinity_flat_line_flag:standard_name = "sea_water_salinity status_flag" ;
	byte qartod_salinity_rate_of_change_flag(time) ;
		qartod_salinity_rate_of_change_flag:_FillValue = 9b ;
		qartod_salinity_rate_of_change_flag:long_name = "QARTOD salinity rate of change test" ;
		qartod_salinity_rate_of_change_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_salinity_rate_of_change_flag:valid_min = 1b ;
		qartod_salinity_rate_of_change_flag:valid_max = 4b ;
		qartod_salinity_rate_of_change_flag:flag_values = 1b, 3b, 4b ;
		qartod_salinity_rate_of_change_flag:comment = "QARTOD salinity rate of change test" ;
		qartod_salinity_rate_of_change_flag:standard_name = "sea_water_salinity status_flag" ;
	byte qartod_salinity_spike_flag(time) ;
		qartod_salinity_spike_flag:_FillValue = 9b ;
		qartod_salinity_spike_flag:long_name = "QARTOD salinity spike test" ;
		qartod_salinity_spike_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_salinity_spike_flag:valid_min = 1b ;
		qartod_salinity_spike_flag:valid_max = 4b ;
		qartod_salinity_spike_flag:flag_values = 1b, 3b, 4b ;
		qartod_salinity_spike_flag:comment = "QARTOD salinity spike test" ;
		qartod_salinity_spike_flag:standard_name = "sea_water_salinity status_flag" ;
	byte qartod_syntax_flag ;
		qartod_syntax_flag:_FillValue = 9b ;
		qartod_syntax_flag:long_name = "QARTOD syntax test" ;
		qartod_syntax_flag:flag_meanings = "Pass Fail" ;
		qartod_syntax_flag:valid_min = 1b ;
		qartod_syntax_flag:valid_max = 4b ;
		qartod_syntax_flag:flag_values = 1b, 4b ;
		qartod_syntax_flag:comment = "QARTOD syntax test" ;
	byte qartod_temperature_climatological_flag(time) ;
		qartod_temperature_climatological_flag:_FillValue = 9b ;
		qartod_temperature_climatological_flag:long_name = "QARTOD temperature climatological test" ;
		qartod_temperature_climatological_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_temperature_climatological_flag:valid_min = 1b ;
		qartod_temperature_climatological_flag:valid_max = 4b ;
		qartod_temperature_climatological_flag:flag_values = 1b, 3b, 4b ;
		qartod_temperature_climatological_flag:comment = "QARTOD temperature climatological test" ;
		qartod_temperature_climatological_flag:standard_name = "sea_water_temperature status_flag" ;
	byte qartod_temperature_flat_line_flag(time) ;
		qartod_temperature_flat_line_flag:_FillValue = 9b ;
		qartod_temperature_flat_line_flag:long_name = "QARTOD temperature flat line test" ;
		qartod_temperature_flat_line_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_temperature_flat_line_flag:valid_min = 1b ;
		qartod_temperature_flat_line_flag:valid_max = 4b ;
		qartod_temperature_flat_line_flag:flag_values = 1b, 3b, 4b ;
		qartod_temperature_flat_line_flag:comment = "QARTOD temperature flat line test" ;
		qartod_temperature_flat_line_flag:standard_name = "sea_water_temperature status_flag" ;
	byte qartod_temperature_gross_range_flag(time) ;
		qartod_temperature_gross_range_flag:_FillValue = 9b ;
		qartod_temperature_gross_range_flag:long_name = "QARTOD temperature gross range test" ;
		qartod_temperature_gross_range_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_temperature_gross_range_flag:valid_min = 1b ;
		qartod_temperature_gross_range_flag:valid_max = 4b ;
		qartod_temperature_gross_range_flag:flag_values = 1b, 3b, 4b ;
		qartod_temperature_gross_range_flag:comment = "QARTOD temperature gross range test" ;
		qartod_temperature_gross_range_flag:standard_name = "sea_water_temperature status_flag" ;
	byte qartod_temperature_rate_of_change_flag(time) ;
		qartod_temperature_rate_of_change_flag:_FillValue = 9b ;
		qartod_temperature_rate_of_change_flag:long_name = "QARTOD temperature rate of change test" ;
		qartod_temperature_rate_of_change_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_temperature_rate_of_change_flag:valid_min = 1b ;
		qartod_temperature_rate_of_change_flag:valid_max = 4b ;
		qartod_temperature_rate_of_change_flag:flag_values = 1b, 3b, 4b ;
		qartod_temperature_rate_of_change_flag:comment = "QARTOD temperature rate of change test" ;
		qartod_temperature_rate_of_change_flag:standard_name = "sea_water_temperature status_flag" ;
	byte qartod_temperature_spike_flag(time) ;
		qartod_temperature_spike_flag:_FillValue = 9b ;
		qartod_temperature_spike_flag:long_name = "QARTOD temperature spike test" ;
		qartod_temperature_spike_flag:flag_meanings = "Pass Suspect Fail" ;
		qartod_temperature_spike_flag:valid_min = 1b ;
		qartod_temperature_spike_flag:valid_max = 4b ;
		qartod_temperature_spike_flag:flag_values = 1b, 3b, 4b ;
		qartod_temperature_spike_flag:comment = "QARTOD temperature spike test" ;
		qartod_temperature_spike_flag:standard_name = "sea_water_temperature status_flag" ;
	byte qartod_timing_and_gap_flag ;
		qartod_timing_and_gap_flag:_FillValue = 9b ;
		qartod_timing_and_gap_flag:long_name = "QARTOD timing and gap test" ;
		qartod_timing_and_gap_flag:flag_meanings = "Pass Fail" ;
		qartod_timing_and_gap_flag:valid_min = 1b ;
		qartod_timing_and_gap_flag:valid_max = 4b ;
		qartod_timing_and_gap_flag:flag_values = 1b, 4b ;
		qartod_timing_and_gap_flag:comment = "QARTOD timing and gap test" ;

// global attributes:
		:Conventions = "CF-1.6, Unidata Dataset Discovery v1.0" ;
		:Metadata_Conventions = "CF-1.6, Unidata Dataset Discovery v1.0" ;
		:acknowledgement = "This deployment supported by ..." ;              // Free-text attribution
        :comment = " " ;                                                     // Any additional notes you may have to describe the dataset
        :contributor_name = " " ;                                            // Comma-separated list of contirbutor names
        :contributor_role = " " ;                                            // Comma-separated list of roles for each contributor listed in contributor_names
        :creator_email = " " ;                                               // E-Mail address of the creator responsible for the dataset
        :creator_name = " " ;                                                // Name of the creator
        :creator_url = " " ;                                                 // The URL of the person (or other creator type specified by the creator_type attribute) principally responsible for creating this data. 
        :date_created = " " ;                                                // ISO-8601 Date string for when the dataset was created
		:date_issued = " " ;                                                 // ISO-8601 Date string for when the dataset was issued
		:date_modified = " " ;                                               // ISO-8601 Date string for when the dataset was last modified
        :format_version = "IOOS_Glider_NetCDF_v3.0-qartod" ;
        :history = " " ;                                                     // List of strings describing historical modifications ot the dataset
        :id = " " ;                                                          // GliderDAC Deployment Identifier, e.g. ru29-20150318T0312
        :institution = " " ;                                                 // Institution responsible for this dataset
        :ioos_regional_association = " " ;                                   // IOOS Regional Association that is associated with this dataset
        :keywords = "AUVS > Autonomous Underwater Vehicles, Oceans > Ocean Pressure > Water Pressure, Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Conductivity, Oceans > Salinity/Density > Density, Oceans > Salinity/Density > Salinity" ;
        :keywords_vocabulary = "GCMD Science Keywords" ;
        :license = "This data may be redistributed and used without restriction.  Data provided as is with no expressed or implied assurance of quality assurance or quality control" ; // Provide the URL to a standard or specific license, enter "Freely Distributed" or "None", or describe any restrictions to data access and distribution in free text.
        :metadata_link = "https://github.com/ioos/ioosngdac/" ;              // Link to the Metadata specification for GliderDAC
        :naming_authority = "gov.noaa.ioos" ;                                // The organization that provides the initial id (see above) for the dataset. The naming authority should be uniquely specified by this attribute. We recommend using reverse-DNS naming for the naming authority; URIs are also acceptable. Example: 'edu.ucar.unidata'.
        :platform_type = "Slocum Glider" ;                                   // Type of glider used to make collections
		:processing_level = " " ;
		:project = " " ;                                                     // Project the collection was a part of
		:publisher_email = " " ;                                             // The email address of the person (or other entity specified by the publisher_type attribute) responsible for publishing the data file or product to users, with its current metadata and format.
		:publisher_name = " " ;                                              // The name of the person (or other entity specified by the publisher_type attribute) responsible for publishing the data file or product to users, with its current metadata and format.
		:publisher_url = " " ;                                               // The URL of the person (or other entity specified by the publisher_type attribute) responsible for publishing the data file or product to users, with its current metadata and format.
		:references = "https://ioos.noaa.gov/wp-content/uploads/2015/10/Manual-for-QC-of-Glider-Data_05_09_16.pdf" ;
		:sea_name = " " ;                                                    // The name of the sea in which the data were collected. See https://www.nodc.noaa.gov/General/NODC-Archive/seanamelist.txt for a list of NCEI sea names
		:source = "Observational data from a profiling glider" ;             // The method of production of the original data. If it was model-generated, source should name the model and its version. If it is observational, source should characterize it. This attribute is defined in the CF Conventions. Examples: 'temperature from CTD #1234'; 'world model v.0.1'.
		:standard_name_vocabulary = "CF-v37" ;                               // CF Standard Name table used for this dataset. http://cfconventions.org/documents.html contains a list of table versions.
		:summary = " " ;                                                     // A paragraph describing the dataset, analogous to an abstract for a paper.
		:title = " " ;                                                       // GliderDAC Deployment Identifier
		:wmo_id = " " ;                                                      // WMO Identifier assigned by the WMO office.
}

